* EESchema Netlist Version 1.1 (Spice format) creation date: Sun 10 Feb 2013 02:18:08 PM CET

* To exclude a component from the Spice Netlist add [Spice_Netlist_Enabled] user FIELD set to: N
* To reorder the component spice node sequence add [Spice_Node_Sequence] user FIELD and define sequence: 2,1,0

*Sheet Name:/
C2  6 0 1uF		
C1  6 0 1uF		
P1  6 0 CONN_2		
P3  7 12 8 17 16 14 9 1 CONN_8		
P2  13 10 11 2 15 3 4 18 CONN_8		
XU2  6 15 16 6 3 14 0 9 4 6 1 18 6 6 74LS126		
XU1  6 13 7 6 10 12 0 8 11 6 17 2 6 6 74LS126		

.end
